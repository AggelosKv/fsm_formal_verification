package fsm_stages_pkg;

    typedef enum logic[1:0] { start = 2'b00, odd = 2'b01, even = 2'b10, fin = 2'b11 } c_state; //stages of fsm

endpackage